module ControlHazard(input BranchSel, output Flush);
  assign Flush = BranchSel;
endmodule